module IM(
	A,
	D_out
    );

	input [9:0] A;
	output [31:0] D_out;

	reg [31:0] data [1023:0];	// 256x31 data

	integer i;
	initial begin
		for (i=0;i<1024;i=i+1) data[i] = 'h00000000;
	end
    initial $readmemh("D:/BC.hex", data);
	assign D_out = data[A];

endmodule