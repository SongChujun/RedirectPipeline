`timescale 1ns / 1ns

module controllertb;
    reg[31:0] IR;
    wire[3:0] ALUop;
    wire dmload;
    wire dmstr;
    wire dmsel;
    wire[4:0] ra;
    wire[4:0] rb;
    wire[4:0] rt;
    wire[4:0] rs;
    wire[5:0] funct;
    wire[5:0] op;
    wire[15:0] imm;
    reg clk;
    initial
    begin
     IR<=0;
     IR[31:26]<=6'b110111;
     IR[5:0]<=6'b1001;
     #100
     IR[31:26]<=6'b111111;
     #100
     IR[31:26]<=6'b100011;
     #100
     IR[31:26]<=6'b101011;
    end
    // always@(posedge clk)

//   initial
//    begin
//    IR<=0;
//    #100
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b100000;
//    IR<=0;
//    #100
//    IR[31:26]<=6'b1000;
//    IR<=0;
//    #100
//    IR[31:26]<=6'b1001;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b100001;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b100100;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b1100;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b0;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b11;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b10;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b100010;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b100101;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b1101;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b100111;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b100011;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b101011;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b100;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b101;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b101010;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b1010;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b101011;
//    IR<=0;  
//    #10
//    IR[31:26]<=6'b1010;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b101011;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b10;
//    IR<=0;

//    #10
//    IR[5:0]<=6'b11;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b1000;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b1100;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b0;
//    IR[5:0]<=6'b110;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b1110;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b100100;
//    IR<=0;
//    #10
//    IR[31:26]<=6'b1;
//    IR<=0;
//    end
    always #20 clk <= ~clk;
    controller u1(.IR(IR),.ALUop(ALUop),.dmload(dmload),.dmstr(dmstr),.dmsel(dmsel),.ra(ra),.rb(rb),.rt(rt),.rs(rs),.funct(funct),.op(op),.imm(imm));
endmodule